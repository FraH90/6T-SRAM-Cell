** Profile: "SCHEMATIC1-transient"  [ C:\Users\FraH\Desktop\StorageCircuits\0a-6TCell-SRAM\0a-6tcell-pspicefiles\schematic1\transient.sim ] 

** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\Cadence\LibreriePACE\an35.lib" 
.lib "C:\Cadence\LibreriePACE\ams.lib" 
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
