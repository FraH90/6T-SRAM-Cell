** Profile: "SCHEMATIC1-0a-WriteVerify"  [ C:\Users\FraH\Desktop\StorageCircuits\0b-6TCell-SRAM - RW\0a-6tcell-pspicefiles\schematic1\0a-writeverify.sim ] 

** Creating circuit file "0a-WriteVerify.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\Cadence\LibrerieMatarrese\diodi.lib" 
.lib "C:\Cadence\LibrerieMatarrese\base.lib" 
.lib "C:\Cadence\LibreriePACE\an35.lib" 
.lib "C:\Cadence\LibreriePACE\ams.lib" 
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
